`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:09:00 12/15/2020 
// Design Name: 
// Module Name:    DM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DM(
    input [31:0] A,
    input [31:0] WD,
	 input DMWr,
	 input [31:0] PC,
    input clk,
    input reset,
    output [31:0] D
    );
	reg [31:0] DM[0:4095];
	integer i;
	initial begin
		for(i=0;i<4096;i=i+1) begin
			DM[i] <= 32'b00000000;
		end
	end
	//��ʼ��
	
	always @(posedge clk)begin
		if(reset) begin
			for(i=0;i<4096;i=i+1) begin
				DM[i] <= 32'b0;
			end
		end
		else if(DMWr) begin
			DM[A[13:2]] <= WD;
			$display("%d@%h: *%h <= %h",$time, PC, {A[31:2],2'b00}, WD);
		end
	end
	//DMд�����
	
	assign D = DM[A[13:2]];
endmodule
